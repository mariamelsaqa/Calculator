module final_tb();
reg [8:0] B;
wire [6:0] mux_out;
Final f ();
endmodule
